`include "design.sv"
`include "bitonic_trans.sv"
`include "bitonic_gen.sv"
`include "bitonic_intf.sv"
`include "bitonic_bfm.sv"
`include "bitonic_env.sv"
`include "bitonic_test.sv"
`include "tb_bitonic_tb.sv"





